["Ratione nemo excepturi quis id voluptas dolor. Ipsum necessitatibus sed rerum. Ducimus eum est omnis officiis repellat deserunt beatae.", "Minima qui velit culpa et aliquid. Cupiditate rem nihil adipisci. Sed molestiae nisi placeat non recusandae nemo. Autem ducimus est vel. Excepturi quia fugiat non nam."]